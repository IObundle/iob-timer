//Memory map
`define TIMER_ADDR_W 3
`define TIMER_WDATA_W 1
