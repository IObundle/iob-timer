//Memory map
`define TIMER_ADDR_W 2

`define TIMER_RESET (`TIMER_ADDR_W'd0)
`define TIMER_STOP (`TIMER_ADDR_W'd1)
`define TIMER_DATA_HIGH (`TIMER_ADDR_W'd2)
`define TIMER_DATA_LOW (`TIMER_ADDR_W'd3)

