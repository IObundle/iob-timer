`define TIMER_ADDR_W 2
`define TIMER_WDATA_W 1
`ifndef DATA_W
 `define DATA_W 32
`endif
